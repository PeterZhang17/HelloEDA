rtl need to be added
testbench.sv need to be added
