// Author: Peter
// Version: V0.0.1
// Update on: 01-OCT-2022

module hello;
  initial 
    begin
      $display("Hello, World");
      $finish ;
    end
endmodule
